* R ladder voltage divider
*
* An intentionally simple example which we expect will have
* no states of any kind (differential or algebraic)

.param vdc = 1

V1 in 0 DC 'vdc'
r1 in out 1
r2 out 0 1

.end
